module random_color(
    input logic clock,
    input logic reset,
    output logic [7:0] color 
    );

endmodule