module tb_random_color();
logic clock;
logic reset;
logic [3:0] x;
logic [9:0] rnd;


			
		
	
endmodule
